//*****************************************************************//
// Lookup table for Distributed Arithmetic 
// Created By - Vrishbhan Singh Sisodia
// San Jose State University
// EE 278
//*****************************************************************//
module lut (in_80, out_80);
	input [5:0] in_80;
	output [5:0] out_80;
	wire [5:0] in_80;
	reg [5:0] out_80;
	
	always @(in_80)
	begin
		case (in_80)
			6'b000000: out_80 = 0;
			6'b000001: out_80 = 7;
			6'b000010: out_80 = -7;
			6'b000011: out_80 = 0;
			6'b000100: out_80 = 5;
			6'b000101: out_80 = 12;
			6'b000110: out_80 = -2;
			6'b000111: out_80 = 5;
			6'b001000: out_80 = 5;
			6'b001001: out_80 = 12;
			6'b001010: out_80 = -2;
			6'b001011: out_80 = 5;
			6'b001100: out_80 = 10;
			6'b001101: out_80 = 17;
			6'b001110: out_80 = 3;
			6'b001111: out_80 = 10;
			6'b010000: out_80 = -5;
			6'b010001: out_80 = 2;
			6'b010010: out_80 = -12;
			6'b010011: out_80 = -5;
			6'b010100: out_80 = 0;
			6'b010101: out_80 = 7;
			6'b010110: out_80 = -7;
			6'b010111: out_80 = 0;
			6'b011000: out_80 = 0;
			6'b011001: out_80 = 7;
			6'b011010: out_80 = -7;
			6'b011011: out_80 = 0;
			6'b011100: out_80 = 5;
			6'b011101: out_80 = 12;
			6'b011110: out_80 = -2;
			6'b011111: out_80 = 5;
			6'b100000: out_80 = 3;
			6'b100001: out_80 = 10;
			6'b100010: out_80 = -4;
			6'b100011: out_80 = 3;
			6'b100100: out_80 = 8;
			6'b100101: out_80 = 15;
			6'b100110: out_80 = 1;
			6'b100111: out_80 = 8;
			6'b101000: out_80 = 8;
			6'b101001: out_80 = 15;
			6'b101010: out_80 = 1;
			6'b101011: out_80 = 8;
			6'b101100: out_80 = 13;
			6'b101101: out_80 = 20;
			6'b101110: out_80 = 6;
			6'b101111: out_80 = 13;
			6'b110000: out_80 = -2;
			6'b110001: out_80 = 5;
			6'b110010: out_80 = -9;
			6'b110011: out_80 = -2;
			6'b110100: out_80 = 3;
			6'b110101: out_80 = 10;
			6'b110110: out_80 = -4;
			6'b110111: out_80 = 3;
			6'b111000: out_80 = 3;
			6'b111001: out_80 = 10;
			6'b111010: out_80 = -4;
			6'b111011: out_80 = 3;
			6'b111100: out_80 = 8;
			6'b111101: out_80 = 15;
			6'b111110: out_80 = 1;
			6'b111111: out_80 = 8;
			default: out_80 = 0;
		endcase
	end
endmodule
